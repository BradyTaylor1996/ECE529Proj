SRAM Cell Subcircuit

* Models
.include ./sram_array.txt
.include ./SA_array.txt
.include ./col_devices_array.txt

* Parameters
.param p = 5N
.param dt = 10P

* Voltage Sources
Vpwr vdd gnd 1.8
Vpc pc gnd pwl 0 0 p 0 'p+dt' 1.8 '6*p' 1.8 '6*p+dt' 0 '7*p' 0 '7*p+dt' 1.8 '11*p' 1.8 '11*p+dt' 0 '12*p' 0 '12*p+dt' 1.8 '17*p' 1.8 '17*p+dt' 0 '18*p' 0 '18*p+dt' 1.8
Vw w gnd pwl 0 0 '2*p' 0 '2*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '13*p' 0 '13*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0
Vd0 d0 gnd pwl 0 0 '2*p' 0 '2*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0
Vd1 d1 gnd 0
Vd2 d2 gnd pwl 0 0 '2*p' 0 '2*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0
Vd3 d3 gnd 0
Vd4 d4 gnd pwl 0 0 '2*p' 0 '2*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0
Vd5 d5 gnd 0
Vd6 d6 gnd pwl 0 0 '2*p' 0 '2*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0
Vd7 d7 gnd 0
Vd_bar0 d_bar0 0
Vd_bar1 d_bar1 gnd pwl 0 0 '2*p' 0 '2*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0
Vd_bar2 d_bar2 0
Vd_bar3 d_bar3 gnd pwl 0 0 '2*p' 0 '2*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0
Vd_bar4 d_bar4 0
Vd_bar5 d_bar5 gnd pwl 0 0 '2*p' 0 '2*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0
Vd_bar6 d_bar6 0
Vd_bar7 d_bar7 gnd pwl 0 0 '2*p' 0 '2*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0
Vd33 d33 gnd pwl 0 0 '13*p' 0 '13*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0
Vd34 d34 gnd 0
Vd35 d35 gnd pwl 0 0 '13*p' 0 '13*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0
Vd36 d36 gnd 0
Vd37 d37 gnd pwl 0 0 '13*p' 0 '13*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0
Vd38 d38 gnd 0
Vd39 d39 gnd pwl 0 0 '13*p' 0 '13*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0
Vd40 d40 gnd 0
Vd_bar33 d_bar33 0
Vd_bar34 d_bar34 gnd pwl 0 0 '13*p' 0 '13*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0
Vd_bar35 d_bar35 0
Vd_bar36 d_bar36 gnd pwl 0 0 '13*p' 0 '13*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0
Vd_bar37 d_bar37 0
Vd_bar38 d_bar38 gnd pwl 0 0 '13*p' 0 '13*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0
Vd_bar39 d_bar39 0
Vd_bar40 d_bar40 gnd pwl 0 0 '13*p' 0 '13*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0
Vcol0 col0 gnd pwl 0 0 '3*p' 0 '3*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol1 col1 gnd pwl 0 0 '3*p' 0 '3*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol2 col2 gnd pwl 0 0 '3*p' 0 '3*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol3 col3 gnd pwl 0 0 '3*p' 0 '3*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8 
Vcol4 col4 gnd pwl 0 0 '3*p' 0 '3*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol5 col5 gnd pwl 0 0 '3*p' 0 '3*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol6 col6 gnd pwl 0 0 '3*p' 0 '3*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol7 col7 gnd pwl 0 0 '3*p' 0 '3*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol33 col33 gnd pwl 0 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol34 col34 gnd pwl 0 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol35 col35 gnd pwl 0 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol36 col36 gnd pwl 0 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol37 col37 gnd pwl 0 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol38 col38 gnd pwl 0 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol39 col39 gnd pwl 0 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vcol40 col40 gnd pwl 0 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '14*p' 0 '14*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vsense SenseEnable gnd pwl 0 0 '9*p' 0 '9*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '20*p' 0 '20*p+dt' 1.8
Vwl0 wl0 gnd pwl 0 0 '4*p' 0 '4*p+dt' 1.8 '5*p' 1.8 '5*p+dt' 0 '8*p' 0 '8*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '19*p' 0 '19*p+dt' 1.8
Vwl4 wl4 gnd pwl 0 0 '8*p' 0 '8*p+dt' 1.8 '10*p' 1.8 '10*p+dt' 0 '15*p' 0 '15*p+dt' 1.8 '16*p' 1.8 '16*p+dt' 0 '19*p' 0 '19*p+dt' 1.8
*Vwl wl0 gnd pwl 0 0 500N 0 501N 1.8 1U 1.8 1.001U 0 2U 0
*Vse SenseEnable gnd pwl 0 0 1.5U 0 1.501U 1.8 2U 1.8
*Vse SenseEnable gnd 1.8V

* Initial Conditions
*.ic b0 = 1.8
*.ic b_bar0 = 1.8

* Main Circuit
X1 b255 b254 b253 b252 b251 b250 b249 b248 b247 b246 b245 b244 b243 b242 b241 b240 b239 b238 b237 b236 b235 b234 b233 b232 b231 b230 b229 b228 b227 b226 b225 b224 b223 b222 b221 b220 b219 b218 b217 b216 b215 b214 b213 b212 b211 b210 b209 b208 b207 b206 b205 b204 b203 b202 b201 b200 b199 b198 b197 b196 b195 b194 b193 b192 b191 b190 b189 b188 b187 b186 b185 b184 b183 b182 b181 b180 b179 b178 b177 b176 b175 b174 b173 b172 b171 b170 b169 b168 b167 b166 b165 b164 b163 b162 b161 b160 b159 b158 b157 b156 b155 b154 b153 b152 b151 b150 b149 b148 b147 b146 b145 b144 b143 b142 b141 b140 b139 b138 b137 b136 b135 b134 b133 b132 b131 b130 b129 b128 b127 b126 b125 b124 b123 b122 b121 b120 b119 b118 b117 b116 b115 b114 b113 b112 b111 b110 b109 b108 b107 b106 b105 b104 b103 b102 b101 b100 b99 b98 b97 b96 b95 b94 b93 b92 b91 b90 b89 b88 b87 b86 b85 b84 b83 b82 b81 b80 b79 b78 b77 b76 b75 b74 b73 b72 b71 b70 b69 b68 b67 b66 b65 b64 b63 b62 b61 b60 b59 b58 b57 b56 b55 b54 b53 b52 b51 b50 b49 b48 b47 b46 b45 b44 b43 b42 b41 b40 b39 b38 b37 b36 b35 b34 b33 b32 b31 b30 b29 b28 b27 b26 b25 b24 b23 b22 b21 b20 b19 b18 b17 b16 b15 b14 b13 b12 b11 b10 b9 b8 b7 b6 b5 b4 b3 b2 b1 b0 b_bar255 b_bar254 b_bar253 b_bar252 b_bar251 b_bar250 b_bar249 b_bar248 b_bar247 b_bar246 b_bar245 b_bar244 b_bar243 b_bar242 b_bar241 b_bar240 b_bar239 b_bar238 b_bar237 b_bar236 b_bar235 b_bar234 b_bar233 b_bar232 b_bar231 b_bar230 b_bar229 b_bar228 b_bar227 b_bar226 b_bar225 b_bar224 b_bar223 b_bar222 b_bar221 b_bar220 b_bar219 b_bar218 b_bar217 b_bar216 b_bar215 b_bar214 b_bar213 b_bar212 b_bar211 b_bar210 b_bar209 b_bar208 b_bar207 b_bar206 b_bar205 b_bar204 b_bar203 b_bar202 b_bar201 b_bar200 b_bar199 b_bar198 b_bar197 b_bar196 b_bar195 b_bar194 b_bar193 b_bar192 b_bar191 b_bar190 b_bar189 b_bar188 b_bar187 b_bar186 b_bar185 b_bar184 b_bar183 b_bar182 b_bar181 b_bar180 b_bar179 b_bar178 b_bar177 b_bar176 b_bar175 b_bar174 b_bar173 b_bar172 b_bar171 b_bar170 b_bar169 b_bar168 b_bar167 b_bar166 b_bar165 b_bar164 b_bar163 b_bar162 b_bar161 b_bar160 b_bar159 b_bar158 b_bar157 b_bar156 b_bar155 b_bar154 b_bar153 b_bar152 b_bar151 b_bar150 b_bar149 b_bar148 b_bar147 b_bar146 b_bar145 b_bar144 b_bar143 b_bar142 b_bar141 b_bar140 b_bar139 b_bar138 b_bar137 b_bar136 b_bar135 b_bar134 b_bar133 b_bar132 b_bar131 b_bar130 b_bar129 b_bar128 b_bar127 b_bar126 b_bar125 b_bar124 b_bar123 b_bar122 b_bar121 b_bar120 b_bar119 b_bar118 b_bar117 b_bar116 b_bar115 b_bar114 b_bar113 b_bar112 b_bar111 b_bar110 b_bar109 b_bar108 b_bar107 b_bar106 b_bar105 b_bar104 b_bar103 b_bar102 b_bar101 b_bar100 b_bar99 b_bar98 b_bar97 b_bar96 b_bar95 b_bar94 b_bar93 b_bar92 b_bar91 b_bar90 b_bar89 b_bar88 b_bar87 b_bar86 b_bar85 b_bar84 b_bar83 b_bar82 b_bar81 b_bar80 b_bar79 b_bar78 b_bar77 b_bar76 b_bar75 b_bar74 b_bar73 b_bar72 b_bar71 b_bar70 b_bar69 b_bar68 b_bar67 b_bar66 b_bar65 b_bar64 b_bar63 b_bar62 b_bar61 b_bar60 b_bar59 b_bar58 b_bar57 b_bar56 b_bar55 b_bar54 b_bar53 b_bar52 b_bar51 b_bar50 b_bar49 b_bar48 b_bar47 b_bar46 b_bar45 b_bar44 b_bar43 b_bar42 b_bar41 b_bar40 b_bar39 b_bar38 b_bar37 b_bar36 b_bar35 b_bar34 b_bar33 b_bar32 b_bar31 b_bar30 b_bar29 b_bar28 b_bar27 b_bar26 b_bar25 b_bar24 b_bar23 b_bar22 b_bar21 b_bar20 b_bar19 b_bar18 b_bar17 b_bar16 b_bar15 b_bar14 b_bar13 b_bar12 b_bar11 b_bar10 b_bar9 b_bar8 b_bar7 b_bar6 b_bar5 b_bar4 b_bar3 b_bar2 b_bar1 b_bar0 wl255 wl254 wl253 wl252 wl251 wl250 wl249 wl248 wl247 wl246 wl245 wl244 wl243 wl242 wl241 wl240 wl239 wl238 wl237 wl236 wl235 wl234 wl233 wl232 wl231 wl230 wl229 wl228 wl227 wl226 wl225 wl224 wl223 wl222 wl221 wl220 wl219 wl218 wl217 wl216 wl215 wl214 wl213 wl212 wl211 wl210 wl209 wl208 wl207 wl206 wl205 wl204 wl203 wl202 wl201 wl200 wl199 wl198 wl197 wl196 wl195 wl194 wl193 wl192 wl191 wl190 wl189 wl188 wl187 wl186 wl185 wl184 wl183 wl182 wl181 wl180 wl179 wl178 wl177 wl176 wl175 wl174 wl173 wl172 wl171 wl170 wl169 wl168 wl167 wl166 wl165 wl164 wl163 wl162 wl161 wl160 wl159 wl158 wl157 wl156 wl155 wl154 wl153 wl152 wl151 wl150 wl149 wl148 wl147 wl146 wl145 wl144 wl143 wl142 wl141 wl140 wl139 wl138 wl137 wl136 wl135 wl134 wl133 wl132 wl131 wl130 wl129 wl128 wl127 wl126 wl125 wl124 wl123 wl122 wl121 wl120 wl119 wl118 wl117 wl116 wl115 wl114 wl113 wl112 wl111 wl110 wl109 wl108 wl107 wl106 wl105 wl104 wl103 wl102 wl101 wl100 wl99 wl98 wl97 wl96 wl95 wl94 wl93 wl92 wl91 wl90 wl89 wl88 wl87 wl86 wl85 wl84 wl83 wl82 wl81 wl80 wl79 wl78 wl77 wl76 wl75 wl74 wl73 wl72 wl71 wl70 wl69 wl68 wl67 wl66 wl65 wl64 wl63 wl62 wl61 wl60 wl59 wl58 wl57 wl56 wl55 wl54 wl53 wl52 wl51 wl50 wl49 wl48 wl47 wl46 wl45 wl44 wl43 wl42 wl41 wl40 wl39 wl38 wl37 wl36 wl35 wl34 wl33 wl32 wl31 wl30 wl29 wl28 wl27 wl26 wl25 wl24 wl23 wl22 wl21 wl20 wl19 wl18 wl17 wl16 wl15 wl14 wl13 wl12 wl11 wl10 wl9 wl8 wl7 wl6 wl5 wl4 wl3 wl2 wl1 wl0 vdd gnd sram_array

*X2 b b_bar Sense Sense_bar SenseEnable vdd gnd SA_l

X2 b255 b254 b253 b252 b251 b250 b249 b248 b247 b246 b245 b244 b243 b242 b241 b240 b239 b238 b237 b236 b235 b234 b233 b232 b231 b230 b229 b228 b227 b226 b225 b224 b223 b222 b221 b220 b219 b218 b217 b216 b215 b214 b213 b212 b211 b210 b209 b208 b207 b206 b205 b204 b203 b202 b201 b200 b199 b198 b197 b196 b195 b194 b193 b192 b191 b190 b189 b188 b187 b186 b185 b184 b183 b182 b181 b180 b179 b178 b177 b176 b175 b174 b173 b172 b171 b170 b169 b168 b167 b166 b165 b164 b163 b162 b161 b160 b159 b158 b157 b156 b155 b154 b153 b152 b151 b150 b149 b148 b147 b146 b145 b144 b143 b142 b141 b140 b139 b138 b137 b136 b135 b134 b133 b132 b131 b130 b129 b128 b127 b126 b125 b124 b123 b122 b121 b120 b119 b118 b117 b116 b115 b114 b113 b112 b111 b110 b109 b108 b107 b106 b105 b104 b103 b102 b101 b100 b99 b98 b97 b96 b95 b94 b93 b92 b91 b90 b89 b88 b87 b86 b85 b84 b83 b82 b81 b80 b79 b78 b77 b76 b75 b74 b73 b72 b71 b70 b69 b68 b67 b66 b65 b64 b63 b62 b61 b60 b59 b58 b57 b56 b55 b54 b53 b52 b51 b50 b49 b48 b47 b46 b45 b44 b43 b42 b41 b40 b39 b38 b37 b36 b35 b34 b33 b32 b31 b30 b29 b28 b27 b26 b25 b24 b23 b22 b21 b20 b19 b18 b17 b16 b15 b14 b13 b12 b11 b10 b9 b8 b7 b6 b5 b4 b3 b2 b1 b0 b_bar255 b_bar254 b_bar253 b_bar252 b_bar251 b_bar250 b_bar249 b_bar248 b_bar247 b_bar246 b_bar245 b_bar244 b_bar243 b_bar242 b_bar241 b_bar240 b_bar239 b_bar238 b_bar237 b_bar236 b_bar235 b_bar234 b_bar233 b_bar232 b_bar231 b_bar230 b_bar229 b_bar228 b_bar227 b_bar226 b_bar225 b_bar224 b_bar223 b_bar222 b_bar221 b_bar220 b_bar219 b_bar218 b_bar217 b_bar216 b_bar215 b_bar214 b_bar213 b_bar212 b_bar211 b_bar210 b_bar209 b_bar208 b_bar207 b_bar206 b_bar205 b_bar204 b_bar203 b_bar202 b_bar201 b_bar200 b_bar199 b_bar198 b_bar197 b_bar196 b_bar195 b_bar194 b_bar193 b_bar192 b_bar191 b_bar190 b_bar189 b_bar188 b_bar187 b_bar186 b_bar185 b_bar184 b_bar183 b_bar182 b_bar181 b_bar180 b_bar179 b_bar178 b_bar177 b_bar176 b_bar175 b_bar174 b_bar173 b_bar172 b_bar171 b_bar170 b_bar169 b_bar168 b_bar167 b_bar166 b_bar165 b_bar164 b_bar163 b_bar162 b_bar161 b_bar160 b_bar159 b_bar158 b_bar157 b_bar156 b_bar155 b_bar154 b_bar153 b_bar152 b_bar151 b_bar150 b_bar149 b_bar148 b_bar147 b_bar146 b_bar145 b_bar144 b_bar143 b_bar142 b_bar141 b_bar140 b_bar139 b_bar138 b_bar137 b_bar136 b_bar135 b_bar134 b_bar133 b_bar132 b_bar131 b_bar130 b_bar129 b_bar128 b_bar127 b_bar126 b_bar125 b_bar124 b_bar123 b_bar122 b_bar121 b_bar120 b_bar119 b_bar118 b_bar117 b_bar116 b_bar115 b_bar114 b_bar113 b_bar112 b_bar111 b_bar110 b_bar109 b_bar108 b_bar107 b_bar106 b_bar105 b_bar104 b_bar103 b_bar102 b_bar101 b_bar100 b_bar99 b_bar98 b_bar97 b_bar96 b_bar95 b_bar94 b_bar93 b_bar92 b_bar91 b_bar90 b_bar89 b_bar88 b_bar87 b_bar86 b_bar85 b_bar84 b_bar83 b_bar82 b_bar81 b_bar80 b_bar79 b_bar78 b_bar77 b_bar76 b_bar75 b_bar74 b_bar73 b_bar72 b_bar71 b_bar70 b_bar69 b_bar68 b_bar67 b_bar66 b_bar65 b_bar64 b_bar63 b_bar62 b_bar61 b_bar60 b_bar59 b_bar58 b_bar57 b_bar56 b_bar55 b_bar54 b_bar53 b_bar52 b_bar51 b_bar50 b_bar49 b_bar48 b_bar47 b_bar46 b_bar45 b_bar44 b_bar43 b_bar42 b_bar41 b_bar40 b_bar39 b_bar38 b_bar37 b_bar36 b_bar35 b_bar34 b_bar33 b_bar32 b_bar31 b_bar30 b_bar29 b_bar28 b_bar27 b_bar26 b_bar25 b_bar24 b_bar23 b_bar22 b_bar21 b_bar20 b_bar19 b_bar18 b_bar17 b_bar16 b_bar15 b_bar14 b_bar13 b_bar12 b_bar11 b_bar10 b_bar9 b_bar8 b_bar7 b_bar6 b_bar5 b_bar4 b_bar3 b_bar2 b_bar1 b_bar0 out255 out254 out253 out252 out251 out250 out249 out248 out247 out246 out245 out244 out243 out242 out241 out240 out239 out238 out237 out236 out235 out234 out233 out232 out231 out230 out229 out228 out227 out226 out225 out224 out223 out222 out221 out220 out219 out218 out217 out216 out215 out214 out213 out212 out211 out210 out209 out208 out207 out206 out205 out204 out203 out202 out201 out200 out199 out198 out197 out196 out195 out194 out193 out192 out191 out190 out189 out188 out187 out186 out185 out184 out183 out182 out181 out180 out179 out178 out177 out176 out175 out174 out173 out172 out171 out170 out169 out168 out167 out166 out165 out164 out163 out162 out161 out160 out159 out158 out157 out156 out155 out154 out153 out152 out151 out150 out149 out148 out147 out146 out145 out144 out143 out142 out141 out140 out139 out138 out137 out136 out135 out134 out133 out132 out131 out130 out129 out128 out127 out126 out125 out124 out123 out122 out121 out120 out119 out118 out117 out116 out115 out114 out113 out112 out111 out110 out109 out108 out107 out106 out105 out104 out103 out102 out101 out100 out99 out98 out97 out96 out95 out94 out93 out92 out91 out90 out89 out88 out87 out86 out85 out84 out83 out82 out81 out80 out79 out78 out77 out76 out75 out74 out73 out72 out71 out70 out69 out68 out67 out66 out65 out64 out63 out62 out61 out60 out59 out58 out57 out56 out55 out54 out53 out52 out51 out50 out49 out48 out47 out46 out45 out44 out43 out42 out41 out40 out39 out38 out37 out36 out35 out34 out33 out32 out31 out30 out29 out28 out27 out26 out25 out24 out23 out22 out21 out20 out19 out18 out17 out16 out15 out14 out13 out12 out11 out10 out9 out8 out7 out6 out5 out4 out3 out2 out1 out0 SenseEnable vdd gnd SA_array

X3 col255 col254 col253 col252 col251 col250 col249 col248 col247 col246 col245 col244 col243 col242 col241 col240 col239 col238 col237 col236 col235 col234 col233 col232 col231 col230 col229 col228 col227 col226 col225 col224 col223 col222 col221 col220 col219 col218 col217 col216 col215 col214 col213 col212 col211 col210 col209 col208 col207 col206 col205 col204 col203 col202 col201 col200 col199 col198 col197 col196 col195 col194 col193 col192 col191 col190 col189 col188 col187 col186 col185 col184 col183 col182 col181 col180 col179 col178 col177 col176 col175 col174 col173 col172 col171 col170 col169 col168 col167 col166 col165 col164 col163 col162 col161 col160 col159 col158 col157 col156 col155 col154 col153 col152 col151 col150 col149 col148 col147 col146 col145 col144 col143 col142 col141 col140 col139 col138 col137 col136 col135 col134 col133 col132 col131 col130 col129 col128 col127 col126 col125 col124 col123 col122 col121 col120 col119 col118 col117 col116 col115 col114 col113 col112 col111 col110 col109 col108 col107 col106 col105 col104 col103 col102 col101 col100 col99 col98 col97 col96 col95 col94 col93 col92 col91 col90 col89 col88 col87 col86 col85 col84 col83 col82 col81 col80 col79 col78 col77 col76 col75 col74 col73 col72 col71 col70 col69 col68 col67 col66 col65 col64 col63 col62 col61 col60 col59 col58 col57 col56 col55 col54 col53 col52 col51 col50 col49 col48 col47 col46 col45 col44 col43 col42 col41 col40 col39 col38 col37 col36 col35 col34 col33 col32 col31 col30 col29 col28 col27 col26 col25 col24 col23 col22 col21 col20 col19 col18 col17 col16 col15 col14 col13 col12 col11 col10 col9 col8 col7 col6 col5 col4 col3 col2 col1 col0 w d255 d254 d253 d252 d251 d250 d249 d248 d247 d246 d245 d244 d243 d242 d241 d240 d239 d238 d237 d236 d235 d234 d233 d232 d231 d230 d229 d228 d227 d226 d225 d224 d223 d222 d221 d220 d219 d218 d217 d216 d215 d214 d213 d212 d211 d210 d209 d208 d207 d206 d205 d204 d203 d202 d201 d200 d199 d198 d197 d196 d195 d194 d193 d192 d191 d190 d189 d188 d187 d186 d185 d184 d183 d182 d181 d180 d179 d178 d177 d176 d175 d174 d173 d172 d171 d170 d169 d168 d167 d166 d165 d164 d163 d162 d161 d160 d159 d158 d157 d156 d155 d154 d153 d152 d151 d150 d149 d148 d147 d146 d145 d144 d143 d142 d141 d140 d139 d138 d137 d136 d135 d134 d133 d132 d131 d130 d129 d128 d127 d126 d125 d124 d123 d122 d121 d120 d119 d118 d117 d116 d115 d114 d113 d112 d111 d110 d109 d108 d107 d106 d105 d104 d103 d102 d101 d100 d99 d98 d97 d96 d95 d94 d93 d92 d91 d90 d89 d88 d87 d86 d85 d84 d83 d82 d81 d80 d79 d78 d77 d76 d75 d74 d73 d72 d71 d70 d69 d68 d67 d66 d65 d64 d63 d62 d61 d60 d59 d58 d57 d56 d55 d54 d53 d52 d51 d50 d49 d48 d47 d46 d45 d44 d43 d42 d41 d40 d39 d38 d37 d36 d35 d34 d33 d32 d31 d30 d29 d28 d27 d26 d25 d24 d23 d22 d21 d20 d19 d18 d17 d16 d15 d14 d13 d12 d11 d10 d9 d8 d7 d6 d5 d4 d3 d2 d1 d0 d_bar255 d_bar254 d_bar253 d_bar252 d_bar251 d_bar250 d_bar249 d_bar248 d_bar247 d_bar246 d_bar245 d_bar244 d_bar243 d_bar242 d_bar241 d_bar240 d_bar239 d_bar238 d_bar237 d_bar236 d_bar235 d_bar234 d_bar233 d_bar232 d_bar231 d_bar230 d_bar229 d_bar228 d_bar227 d_bar226 d_bar225 d_bar224 d_bar223 d_bar222 d_bar221 d_bar220 d_bar219 d_bar218 d_bar217 d_bar216 d_bar215 d_bar214 d_bar213 d_bar212 d_bar211 d_bar210 d_bar209 d_bar208 d_bar207 d_bar206 d_bar205 d_bar204 d_bar203 d_bar202 d_bar201 d_bar200 d_bar199 d_bar198 d_bar197 d_bar196 d_bar195 d_bar194 d_bar193 d_bar192 d_bar191 d_bar190 d_bar189 d_bar188 d_bar187 d_bar186 d_bar185 d_bar184 d_bar183 d_bar182 d_bar181 d_bar180 d_bar179 d_bar178 d_bar177 d_bar176 d_bar175 d_bar174 d_bar173 d_bar172 d_bar171 d_bar170 d_bar169 d_bar168 d_bar167 d_bar166 d_bar165 d_bar164 d_bar163 d_bar162 d_bar161 d_bar160 d_bar159 d_bar158 d_bar157 d_bar156 d_bar155 d_bar154 d_bar153 d_bar152 d_bar151 d_bar150 d_bar149 d_bar148 d_bar147 d_bar146 d_bar145 d_bar144 d_bar143 d_bar142 d_bar141 d_bar140 d_bar139 d_bar138 d_bar137 d_bar136 d_bar135 d_bar134 d_bar133 d_bar132 d_bar131 d_bar130 d_bar129 d_bar128 d_bar127 d_bar126 d_bar125 d_bar124 d_bar123 d_bar122 d_bar121 d_bar120 d_bar119 d_bar118 d_bar117 d_bar116 d_bar115 d_bar114 d_bar113 d_bar112 d_bar111 d_bar110 d_bar109 d_bar108 d_bar107 d_bar106 d_bar105 d_bar104 d_bar103 d_bar102 d_bar101 d_bar100 d_bar99 d_bar98 d_bar97 d_bar96 d_bar95 d_bar94 d_bar93 d_bar92 d_bar91 d_bar90 d_bar89 d_bar88 d_bar87 d_bar86 d_bar85 d_bar84 d_bar83 d_bar82 d_bar81 d_bar80 d_bar79 d_bar78 d_bar77 d_bar76 d_bar75 d_bar74 d_bar73 d_bar72 d_bar71 d_bar70 d_bar69 d_bar68 d_bar67 d_bar66 d_bar65 d_bar64 d_bar63 d_bar62 d_bar61 d_bar60 d_bar59 d_bar58 d_bar57 d_bar56 d_bar55 d_bar54 d_bar53 d_bar52 d_bar51 d_bar50 d_bar49 d_bar48 d_bar47 d_bar46 d_bar45 d_bar44 d_bar43 d_bar42 d_bar41 d_bar40 d_bar39 d_bar38 d_bar37 d_bar36 d_bar35 d_bar34 d_bar33 d_bar32 d_bar31 d_bar30 d_bar29 d_bar28 d_bar27 d_bar26 d_bar25 d_bar24 d_bar23 d_bar22 d_bar21 d_bar20 d_bar19 d_bar18 d_bar17 d_bar16 d_bar15 d_bar14 d_bar13 d_bar12 d_bar11 d_bar10 d_bar9 d_bar8 d_bar7 d_bar6 d_bar5 d_bar4 d_bar3 d_bar2 d_bar1 d_bar0 b255 b254 b253 b252 b251 b250 b249 b248 b247 b246 b245 b244 b243 b242 b241 b240 b239 b238 b237 b236 b235 b234 b233 b232 b231 b230 b229 b228 b227 b226 b225 b224 b223 b222 b221 b220 b219 b218 b217 b216 b215 b214 b213 b212 b211 b210 b209 b208 b207 b206 b205 b204 b203 b202 b201 b200 b199 b198 b197 b196 b195 b194 b193 b192 b191 b190 b189 b188 b187 b186 b185 b184 b183 b182 b181 b180 b179 b178 b177 b176 b175 b174 b173 b172 b171 b170 b169 b168 b167 b166 b165 b164 b163 b162 b161 b160 b159 b158 b157 b156 b155 b154 b153 b152 b151 b150 b149 b148 b147 b146 b145 b144 b143 b142 b141 b140 b139 b138 b137 b136 b135 b134 b133 b132 b131 b130 b129 b128 b127 b126 b125 b124 b123 b122 b121 b120 b119 b118 b117 b116 b115 b114 b113 b112 b111 b110 b109 b108 b107 b106 b105 b104 b103 b102 b101 b100 b99 b98 b97 b96 b95 b94 b93 b92 b91 b90 b89 b88 b87 b86 b85 b84 b83 b82 b81 b80 b79 b78 b77 b76 b75 b74 b73 b72 b71 b70 b69 b68 b67 b66 b65 b64 b63 b62 b61 b60 b59 b58 b57 b56 b55 b54 b53 b52 b51 b50 b49 b48 b47 b46 b45 b44 b43 b42 b41 b40 b39 b38 b37 b36 b35 b34 b33 b32 b31 b30 b29 b28 b27 b26 b25 b24 b23 b22 b21 b20 b19 b18 b17 b16 b15 b14 b13 b12 b11 b10 b9 b8 b7 b6 b5 b4 b3 b2 b1 b0 b_bar255 b_bar254 b_bar253 b_bar252 b_bar251 b_bar250 b_bar249 b_bar248 b_bar247 b_bar246 b_bar245 b_bar244 b_bar243 b_bar242 b_bar241 b_bar240 b_bar239 b_bar238 b_bar237 b_bar236 b_bar235 b_bar234 b_bar233 b_bar232 b_bar231 b_bar230 b_bar229 b_bar228 b_bar227 b_bar226 b_bar225 b_bar224 b_bar223 b_bar222 b_bar221 b_bar220 b_bar219 b_bar218 b_bar217 b_bar216 b_bar215 b_bar214 b_bar213 b_bar212 b_bar211 b_bar210 b_bar209 b_bar208 b_bar207 b_bar206 b_bar205 b_bar204 b_bar203 b_bar202 b_bar201 b_bar200 b_bar199 b_bar198 b_bar197 b_bar196 b_bar195 b_bar194 b_bar193 b_bar192 b_bar191 b_bar190 b_bar189 b_bar188 b_bar187 b_bar186 b_bar185 b_bar184 b_bar183 b_bar182 b_bar181 b_bar180 b_bar179 b_bar178 b_bar177 b_bar176 b_bar175 b_bar174 b_bar173 b_bar172 b_bar171 b_bar170 b_bar169 b_bar168 b_bar167 b_bar166 b_bar165 b_bar164 b_bar163 b_bar162 b_bar161 b_bar160 b_bar159 b_bar158 b_bar157 b_bar156 b_bar155 b_bar154 b_bar153 b_bar152 b_bar151 b_bar150 b_bar149 b_bar148 b_bar147 b_bar146 b_bar145 b_bar144 b_bar143 b_bar142 b_bar141 b_bar140 b_bar139 b_bar138 b_bar137 b_bar136 b_bar135 b_bar134 b_bar133 b_bar132 b_bar131 b_bar130 b_bar129 b_bar128 b_bar127 b_bar126 b_bar125 b_bar124 b_bar123 b_bar122 b_bar121 b_bar120 b_bar119 b_bar118 b_bar117 b_bar116 b_bar115 b_bar114 b_bar113 b_bar112 b_bar111 b_bar110 b_bar109 b_bar108 b_bar107 b_bar106 b_bar105 b_bar104 b_bar103 b_bar102 b_bar101 b_bar100 b_bar99 b_bar98 b_bar97 b_bar96 b_bar95 b_bar94 b_bar93 b_bar92 b_bar91 b_bar90 b_bar89 b_bar88 b_bar87 b_bar86 b_bar85 b_bar84 b_bar83 b_bar82 b_bar81 b_bar80 b_bar79 b_bar78 b_bar77 b_bar76 b_bar75 b_bar74 b_bar73 b_bar72 b_bar71 b_bar70 b_bar69 b_bar68 b_bar67 b_bar66 b_bar65 b_bar64 b_bar63 b_bar62 b_bar61 b_bar60 b_bar59 b_bar58 b_bar57 b_bar56 b_bar55 b_bar54 b_bar53 b_bar52 b_bar51 b_bar50 b_bar49 b_bar48 b_bar47 b_bar46 b_bar45 b_bar44 b_bar43 b_bar42 b_bar41 b_bar40 b_bar39 b_bar38 b_bar37 b_bar36 b_bar35 b_bar34 b_bar33 b_bar32 b_bar31 b_bar30 b_bar29 b_bar28 b_bar27 b_bar26 b_bar25 b_bar24 b_bar23 b_bar22 b_bar21 b_bar20 b_bar19 b_bar18 b_bar17 b_bar16 b_bar15 b_bar14 b_bar13 b_bar12 b_bar11 b_bar10 b_bar9 b_bar8 b_bar7 b_bar6 b_bar5 b_bar4 b_bar3 b_bar2 b_bar1 b_bar0 vdd gnd WD_array

X4 pc b255 b254 b253 b252 b251 b250 b249 b248 b247 b246 b245 b244 b243 b242 b241 b240 b239 b238 b237 b236 b235 b234 b233 b232 b231 b230 b229 b228 b227 b226 b225 b224 b223 b222 b221 b220 b219 b218 b217 b216 b215 b214 b213 b212 b211 b210 b209 b208 b207 b206 b205 b204 b203 b202 b201 b200 b199 b198 b197 b196 b195 b194 b193 b192 b191 b190 b189 b188 b187 b186 b185 b184 b183 b182 b181 b180 b179 b178 b177 b176 b175 b174 b173 b172 b171 b170 b169 b168 b167 b166 b165 b164 b163 b162 b161 b160 b159 b158 b157 b156 b155 b154 b153 b152 b151 b150 b149 b148 b147 b146 b145 b144 b143 b142 b141 b140 b139 b138 b137 b136 b135 b134 b133 b132 b131 b130 b129 b128 b127 b126 b125 b124 b123 b122 b121 b120 b119 b118 b117 b116 b115 b114 b113 b112 b111 b110 b109 b108 b107 b106 b105 b104 b103 b102 b101 b100 b99 b98 b97 b96 b95 b94 b93 b92 b91 b90 b89 b88 b87 b86 b85 b84 b83 b82 b81 b80 b79 b78 b77 b76 b75 b74 b73 b72 b71 b70 b69 b68 b67 b66 b65 b64 b63 b62 b61 b60 b59 b58 b57 b56 b55 b54 b53 b52 b51 b50 b49 b48 b47 b46 b45 b44 b43 b42 b41 b40 b39 b38 b37 b36 b35 b34 b33 b32 b31 b30 b29 b28 b27 b26 b25 b24 b23 b22 b21 b20 b19 b18 b17 b16 b15 b14 b13 b12 b11 b10 b9 b8 b7 b6 b5 b4 b3 b2 b1 b0 b_bar255 b_bar254 b_bar253 b_bar252 b_bar251 b_bar250 b_bar249 b_bar248 b_bar247 b_bar246 b_bar245 b_bar244 b_bar243 b_bar242 b_bar241 b_bar240 b_bar239 b_bar238 b_bar237 b_bar236 b_bar235 b_bar234 b_bar233 b_bar232 b_bar231 b_bar230 b_bar229 b_bar228 b_bar227 b_bar226 b_bar225 b_bar224 b_bar223 b_bar222 b_bar221 b_bar220 b_bar219 b_bar218 b_bar217 b_bar216 b_bar215 b_bar214 b_bar213 b_bar212 b_bar211 b_bar210 b_bar209 b_bar208 b_bar207 b_bar206 b_bar205 b_bar204 b_bar203 b_bar202 b_bar201 b_bar200 b_bar199 b_bar198 b_bar197 b_bar196 b_bar195 b_bar194 b_bar193 b_bar192 b_bar191 b_bar190 b_bar189 b_bar188 b_bar187 b_bar186 b_bar185 b_bar184 b_bar183 b_bar182 b_bar181 b_bar180 b_bar179 b_bar178 b_bar177 b_bar176 b_bar175 b_bar174 b_bar173 b_bar172 b_bar171 b_bar170 b_bar169 b_bar168 b_bar167 b_bar166 b_bar165 b_bar164 b_bar163 b_bar162 b_bar161 b_bar160 b_bar159 b_bar158 b_bar157 b_bar156 b_bar155 b_bar154 b_bar153 b_bar152 b_bar151 b_bar150 b_bar149 b_bar148 b_bar147 b_bar146 b_bar145 b_bar144 b_bar143 b_bar142 b_bar141 b_bar140 b_bar139 b_bar138 b_bar137 b_bar136 b_bar135 b_bar134 b_bar133 b_bar132 b_bar131 b_bar130 b_bar129 b_bar128 b_bar127 b_bar126 b_bar125 b_bar124 b_bar123 b_bar122 b_bar121 b_bar120 b_bar119 b_bar118 b_bar117 b_bar116 b_bar115 b_bar114 b_bar113 b_bar112 b_bar111 b_bar110 b_bar109 b_bar108 b_bar107 b_bar106 b_bar105 b_bar104 b_bar103 b_bar102 b_bar101 b_bar100 b_bar99 b_bar98 b_bar97 b_bar96 b_bar95 b_bar94 b_bar93 b_bar92 b_bar91 b_bar90 b_bar89 b_bar88 b_bar87 b_bar86 b_bar85 b_bar84 b_bar83 b_bar82 b_bar81 b_bar80 b_bar79 b_bar78 b_bar77 b_bar76 b_bar75 b_bar74 b_bar73 b_bar72 b_bar71 b_bar70 b_bar69 b_bar68 b_bar67 b_bar66 b_bar65 b_bar64 b_bar63 b_bar62 b_bar61 b_bar60 b_bar59 b_bar58 b_bar57 b_bar56 b_bar55 b_bar54 b_bar53 b_bar52 b_bar51 b_bar50 b_bar49 b_bar48 b_bar47 b_bar46 b_bar45 b_bar44 b_bar43 b_bar42 b_bar41 b_bar40 b_bar39 b_bar38 b_bar37 b_bar36 b_bar35 b_bar34 b_bar33 b_bar32 b_bar31 b_bar30 b_bar29 b_bar28 b_bar27 b_bar26 b_bar25 b_bar24 b_bar23 b_bar22 b_bar21 b_bar20 b_bar19 b_bar18 b_bar17 b_bar16 b_bar15 b_bar14 b_bar13 b_bar12 b_bar11 b_bar10 b_bar9 b_bar8 b_bar7 b_bar6 b_bar5 b_bar4 b_bar3 b_bar2 b_bar1 b_bar0 vdd gnd PC_array

* Control Options
.options post probe

* Analysis
.tran 10P '22*p'

* Output
.probe tran v(out0) v(out1) v(out2) v(out3) v(out4) v(out5) v(out6) v(out7) v(out33) v(out34) v(out35) v(out36) v(out37) v(out38) v(out39) v(out40) v(pc) v(wl0) v(wl4) v(w) v(SenseEnable) v(d0) v(d1) v(d2) v(d3) v(d4) v(d5) v(d6) v(d7) v(d33) v(d34) v(d35) v(d36) v(d37) v(d38) v(d39) v(d40) v(d_bar0) v(d_bar1) v(d_bar2) v(d_bar3) v(d_bar4) v(d_bar5) v(d_bar6) v(d_bar7) v(d_bar33) v(d_bar34) v(d_bar35) v(d_bar36) v(d_bar37) v(d_bar38) v(d_bar39) v(d_bar40) v(col0) v(col1) v(col2) v(col3) v(col4) v(col5) v(col6) v(col7) v(col33) v(col34) v(col35) v(col36) v(col37) v(col38) v(col39) v(col40)

.end
